--TEMPORARY PLACEHOLDER FOR VHDL CODE
---lab3 project summary
-- inputs:
--		clk 50mhz in
--		mux para seletor de duty cycle
--
--	interno:
--		divisor de frequência (50mhz papra 1hz)
--		funçao para output 7 segmentos
--
--	outputs:
--		dois 7seg (dezena, unidade)
--		1 LED que pisca a cada 5 pulsos de 1hz
--		onda quadrada de 1hz com duty cycle selecionado pelo mux inicial
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity lab3 is
Port ( B0,B1,B2,B3 : in STD_LOGIC;
A,B,C,D,E,F,G : out STD_LOGIC;
CLK : in STD_LOGIC);
end lab3;
 
architecture Behavioral of lab3 is
 
begin

A <= B0 OR B2 OR (B1 AND B3) OR (NOT B1 AND NOT B3);
B <= (NOT B1) OR (NOT B2 AND NOT B3) OR (B2 AND B3);
C <= B1 OR NOT B2 OR B3;
D <= (NOT B1 AND NOT B3) OR (B2 AND NOT B3) OR (B1 AND NOT B2 AND B3) OR (NOT B1 AND B2) OR B0;
E <= (NOT B1 AND NOT B3) OR (B2 AND NOT B3);
F <= B0 OR (NOT B2 AND NOT B3) OR (B1 AND NOT B2) OR (B1 AND NOT B3);
G <= B0 OR (B1 AND NOT B2) OR ( NOT B1 AND B2) OR (B2 AND NOT B3);
 
end Behavioral;
