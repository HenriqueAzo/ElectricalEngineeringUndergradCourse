library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb is end;

architecture testbench of tb is

	component main
    	port (
        A:      in std_logic_vector(3 downto 0);
        B:      in std_logic_vector(3 downto 0);
        Start:  in std_logic;
        Reset:  in std_logic;
        clck:   in std_logic;
        P:      out std_logic_vector(7 downto 0)
        
    );
    end component main;
    
    --declara��o do tempo de clock
    constant PERIODO : time := 10 ns;
    
    --entradas e sa�das tratadas por sinais, na mesma ordem que no componente
    signal sA:   std_logic_vector(3 downto 0);
    signal sB:   std_logic_vector(3 downto 0);
    signal Stt:  std_logic;
    signal Rst:  std_logic;
    signal Clk:  std_logic := '0';
    signal Outp: std_logic_vector(7 downto 0);
    
    begin
    
    --gera��o do clock
    Clk <= not Clk after PERIODO/2;
    
    --assinalando as entradas e sa�das aos sinais tratados
    dut: main port map( 	 A=> sA,
							 B=> sB,
							 Start=> Stt,
							 Reset=> Rst,
                             clck=> Clk,
                             P=> Outp
							);
    
    
    inc: process is
    begin
    wait for 5 ns;
    
    sA <= "0001";
    sB <= "0010";
    Stt<= '1';
    Rst<= '0';
    
    wait for 5 ns;
    
    Stt<= '0';
    
    wait for 200 ns;
    
    report "resultado: " & to_string(Outp);
    
    wait;
    
end process;
end testbench;

